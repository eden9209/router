interface switch_input_if(input logic clock);
    logic [7:0] data_in;
    logic data_status;
    logic reset;
  endinterface