interface switch_output_if(input logic clock);
    logic [7:0] data_out;
    logic ready;
    logic read;
    endinterface