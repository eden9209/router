package switch_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import switch_agent_pkg::*;

  ///include componnet 
  `include "switch_scoreboard.sv"
  `include "switch_env.sv"
  `include "switch_test.sv" 
endpackage